entity clk_led is
port (
signal clock_in : in bit;
signal clock_led : out bit

);
end entity clk_led;


architecture c_clk_led of clk_led is

begin










end architecture c_clk_led;
